module To_7segment (
	input [3:0] data,
  output  [6:0] hex
  );

  assign hex = (data[3:0] == 8'd15) ? 7'b0001110:
              (data[3:0] == 8'd14) ? 7'b0000110:
              (data[3:0] == 8'd13) ? 7'b0100001:
              (data[3:0] == 8'd12) ? 7'b1000110:
              (data[3:0] == 8'd11) ? 7'b0000011:
              (data[3:0] == 8'd10) ? 7'b0001000:
              (data[3:0] == 8'd9) ? 7'b0010000:
              (data[3:0] == 8'd8) ? 7'b0000000:
              (data[3:0] == 8'd7) ? 7'b1111000:
              (data[3:0] == 8'd6) ? 7'b0000010:
              (data[3:0] == 8'd5) ? 7'b0010010:
              (data[3:0] == 8'd4) ? 7'b0011001:
              (data[3:0] == 8'd3) ? 7'b0110000:
              (data[3:0] == 8'd2) ? 7'b0100100:
              (data[3:0] == 8'd1) ? 7'b1111001: 7'b1000000;

endmodule // To_7segmen
