module Instruction_Memory (address,instruction);
input [31:0] address;
output [31:0] instruction;

reg [31:0]mem[0:99];

initial begin
  mem[0]  = 32'b101010_00000_00000_0000000000000011; // JMP $3
  mem[1]  = 32'b000000_00010_00011_00010_00000000000;
  mem[2]  = 32'b100001_00011_00011_0000000000010000;
  mem[3]  = 32'b000001_00101_00011_0000000000010000; // add R5, R3, R0
  mem[4]  = 32'b101010_00000_00000_1111111111111101; // JMP $3
/*
  mem[0]   = 32'b100000_00001_00001_0000000000010000;
  mem[1]   = 32'b000000_00010_00011_00010_00000000000;
  mem[2]   = 32'b100001_00011_00011_0000000000010000;
  mem[3]   = 32'b000001_00101_00011_0000000000010000;
  mem[4]   = 32'b100101_00011_00111_0000000000001001; // store  R3 in M[R7+$9]
  mem[5]   = 32'b100100_00100_00111_0000000000001000; // load  m[15] in r4
  mem[6]   = 32'b101000_00000_00000_0000000000001000; // BEZ R0, R0, $8
  mem[7]   = 32'b101000_00000_00001_0000000000001000; // BEZ R0, R1, $8
  mem[8]   = 32'b101001_00100_00111_0000000000001000; // BNE R4, R7, $8
  mem[9]   = 32'b101001_00100_00100_0000000000001000; // BNE R4, R4, $8
  mem[10]  = 32'b101010_00100_00111_0000000000001000; // JMP $16
  mem[16]  = 32'b101010_00100_00111_0000000000000001; // JMP $1
  */
  /*
  mem[2]  = 32'b000010_00000_00101_00110_00000000000;
  mem[3]  = 32'b000011_00010_00111_01000_00000000000;
  mem[4]  = 32'b000100_00011_01001_01010_00000000000;
  mem[5]  = 32'b000101_00000_01011_01100_00000000000;
  mem[6]  = 32'b000110_00000_01101_01110_00000000000;
  mem[7]  = 32'b000111_00000_01101_01110_00000000000;
  mem[8]  = 32'b001000_00000_01101_01110_00000000000;
  mem[9]  = 32'b001001_00000_01101_01110_00000000000;
  mem[10] = 32'b001010_00000_01101_01110_00000000000;
  mem[11] = 32'b001011_00000_01101_01110_00000000000;
  mem[12] = 32'b001100_00000_01101_01110_00000000000;
  mem[13] = 32'b100000_00000_01101_01110_00000000000;
  mem[14] = 32'b100001_00000_01101_01110_00000000000;
  mem[15] = 32'b100100_00000_01101_01110_00000000000;
  mem[16] = 32'b100101_00000_01101_01110_00000000000;
  mem[17] = 32'b101000_00000_01101_01110_00000000000;
  mem[18] = 32'b101001_00000_01101_01110_00000000000;
  mem[19] = 32'b101010_00000_01101_01110_00000000000;
  
  32'b100000_00001_00000_00000_00000001010;//-- Addi
2. 32'b000001_00010_00000_00001_00000000000;//-- Add
3. 32'b000011_00011_00000_00001_00000000000;//-- sub
4. 32'b000101_00100_00010_00011_00000000000;//-- And
5. 32'b100001_00101_00000_00000_01000110100;//-- Subi
6. 32'b000110_00101_00101_00011_00000000000;//-- or
7. 32'b000111_00110_00101_00000_00000000000;//-- nor
8. 32'b001000_00000_00101_00001_00000000000;//-- xor
9. 32'b001000_00111_00101_00001_00000000000;//-- xor
10. 32'b001001_00111_00100_00010_00000000000;//-- sla
11. 32'b001010_01000_00011_00010_00000000000;//-- sll
12. 32'b001011_01001_00110_00010_00000000000;//-- sra
13. 32'b001100_01010_00110_00010_00000000000;//-- srl
14. 32'b100000_00001_00000_00000_10000000000;//-- Addi
15. 32'b100101_00010_00001_00000_00000000000;//-- st
16. 32'b100100_01011_00001_00000_00000000000;//-- ld
17. 32'b100101_00011_00001_00000_00000000100;//-- st
18. 32'b100101_00100_00001_00000_00000001000;//-- st
19. 32'b100101_00101_00001_00000_00000001100;//-- st
20. 32'b100101_00110_00001_00000_00000010000;//-- st
21. 32'b100101_00111_00001_00000_00000010100;//-- st
22. 32'b100101_01000_00001_00000_00000011000;//-- st
23. 32'b100101_01001_00001_00000_00000011100;//-- st
24. 32'b100101_01010_00001_00000_00000100000;//-- st
25. 32'b100101_01011_00001_00000_00000100100;//-- st
26. 32'b100000_00001_00000_00000_00000000011;//-- Addi
27. 32'b100000_00100_00000_00000_10000000000;//-- Addi
28. 32'b100000_00010_00000_00000_00000000000;//-- Addi
29. 32'b100000_00011_00000_00000_00000000001;//-- Addi
30. 32'b100000_01001_00000_00000_00000000010;//-- Addi
31. 32'b001010_01000_00011_01001_00000000000;//-- sll
32. 32'b000001_01000_00100_01000_00000000000;//-- Add
33. 32'b100100_00101_01000_00000_00000000000;//-- ld
34. 32'b100100_00110_01000_11111_11111111100;//-- ld
35. 32'b000011_01001_00101_00110_00000000000;//-- sub
36. 32'b100000_01010_00000_10000_00000000000;//-- Addi
37. 32'b100000_01011_00000_00000_00000010000;//-- Addi
38. 32'b001010_01010_01010_01011_00000000000;//-- sll
39. 32'b000101_01001_01001_01010_00000000000;//-- And
40. 32'b101000_00000_01001_00000_00000000010;//-- Bez
41. 32'b100101_00101_01000_11111_11111111100;//-- st
  */
  //$readmemb("instruction_file.txt",mem); // readmemh for hex
end

assign instruction = mem[address];

endmodule // InstructionMemorys
